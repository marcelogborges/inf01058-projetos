library verilog;
use verilog.vl_types.all;
entity DIVFREQ_vlg_vec_tst is
end DIVFREQ_vlg_vec_tst;
