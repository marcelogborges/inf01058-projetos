library verilog;
use verilog.vl_types.all;
entity CONTA_A_DOR_vlg_vec_tst is
end CONTA_A_DOR_vlg_vec_tst;
