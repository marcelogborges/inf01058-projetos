library verilog;
use verilog.vl_types.all;
entity LAB03_vlg_vec_tst is
end LAB03_vlg_vec_tst;
