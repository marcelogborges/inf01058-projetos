library verilog;
use verilog.vl_types.all;
entity DIVFREQ_vlg_sample_tst is
    port(
        CLK_IN          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end DIVFREQ_vlg_sample_tst;
